module memory(clk, reset, address, data_in, data_out, read, write, ready);

input clk;
input reset;
input address;
input data_in;
output data_out;
input read;
input write;
output ready;

endmodule
